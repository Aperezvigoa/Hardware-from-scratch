CHIP And {
	IN a, b;
	OUT out;

	PARTS:
	Nand(a= a, b= b, out= aNandb);
	Not(in= aNandb, out= out);
}
