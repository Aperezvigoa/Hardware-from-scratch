CHIP Not {
    IN in;
    OUT out;

    PARTS:
	And(a= in, b= false, out= aAndfalse);
}
